** Profile: "SCHEMATIC1-prelab1"  [ C:\Users\nmunoz\Documents\wsu\EE352\LAB1\PreLab4_ee532-PSpiceFiles\SCHEMATIC1\prelab1.sim ] 

** Creating circuit file "prelab1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\nmunoz\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 1000 1 47.2k
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
